// Copyright lowRISC contributors.
// Copyright 2018 ETH Zurich and University of Bologna, see also CREDITS.md.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`ifdef RISCV_FORMAL
  `define RVFI
`endif

/**
 * Instruction Decode Stage
 *
 * Decode stage of the core. It decodes the instructions and hosts the register
 * file.
 */

`include "prim_assert.sv"
`include "dv_fcov_macros.svh"

module cve2_id_stage #(
  parameter bit               RV32E       = 0,
  parameter cve2_pkg::rv32m_e RV32M       = cve2_pkg::RV32MFast,
  parameter cve2_pkg::rv32b_e RV32B       = cve2_pkg::RV32BNone,
  parameter                   N_HWLP      = 2,
  parameter                   N_HWLP_BITS = $clog2(N_HWLP),
  parameter bit [31:0]        COPROC_OPCODE = 32'h00400400
) (
  input  logic                      clk_i,
  input  logic                      rst_ni,

  input  logic                      fetch_enable_i,
  output logic                      ctrl_busy_o,
  output logic                      illegal_insn_o,

  // Interface to IF stage
  input  logic                      instr_valid_i,
  input  logic [31:0]               instr_rdata_i,         // from IF-ID pipeline registers
  input  logic [31:0]               instr_rdata_alu_i,     // from IF-ID pipeline registers
  input  logic [15:0]               instr_rdata_c_i,       // from IF-ID pipeline registers
  input  logic                      instr_is_compressed_i,
  output logic                      instr_req_o,
  output logic                      instr_first_cycle_id_o,
  output logic                      instr_valid_clear_o,   // kill instr in IF-ID reg
  output logic                      id_in_ready_o,         // ID stage is ready for next instr

  // Jumps and branches
  input  logic                      branch_decision_i,

  // IF and ID stage signals
  output logic                      pc_set_o,
  output cve2_pkg::pc_sel_e         pc_mux_o,
  output cve2_pkg::exc_pc_sel_e     exc_pc_mux_o,
  output cve2_pkg::exc_cause_e      exc_cause_o,

  input  logic                      illegal_c_insn_i,
  input  logic                      instr_fetch_err_i,
  input  logic                      instr_fetch_err_plus2_i,

  input  logic [31:0]               pc_id_i,

  // Stalls
  input  logic                      ex_valid_i,       // EX stage has valid output
  input  logic                      lsu_resp_valid_i, // LSU has valid output, or is done
  // ALU
  output cve2_pkg::alu_op_e         alu_operator_ex_o,
  output logic [31:0]               alu_operand_a_ex_o,
  output logic [31:0]               alu_operand_b_ex_o,



//---------------------------------------------------------------------------------
  output logic [31:0]               alu_operand_c_ex_o,
//---------------------------------------------------------------------------------



  // Multicycle Operation Stage Register
  input  logic [1:0]                imd_val_we_ex_i,
  input  logic [33:0]               imd_val_d_ex_i[2],
  output logic [33:0]               imd_val_q_ex_o[2],

  // MUL, DIV
  output logic                      mult_en_ex_o,
  output logic                      div_en_ex_o,
  output logic                      mult_sel_ex_o,
  output logic                      div_sel_ex_o,
  output cve2_pkg::md_op_e          multdiv_operator_ex_o,
  output logic  [1:0]               multdiv_signed_mode_ex_o,
  output logic [31:0]               multdiv_operand_a_ex_o,
  output logic [31:0]               multdiv_operand_b_ex_o,

  // CSR
  output logic                      csr_access_o,
  output cve2_pkg::csr_op_e         csr_op_o,
  output logic                      csr_op_en_o,
  output logic                      csr_save_if_o,
  output logic                      csr_save_id_o,
  output logic                      csr_restore_mret_id_o,
  output logic                      csr_restore_dret_id_o,
  output logic                      csr_save_cause_o,
  output logic [31:0]               csr_mtval_o,
  input  cve2_pkg::priv_lvl_e       priv_mode_i,
  input  logic                      csr_mstatus_tw_i,
  input  logic                      illegal_csr_insn_i,

  // Interface to load store unit
  output logic                      lsu_req_o,
  output logic                      lsu_we_o,
  output logic [1:0]                lsu_type_o,
  output logic                      lsu_sign_ext_o,
  output logic [31:0]               lsu_wdata_o,



//---------------------------------------------------------------------------------
  //Signals needed for Post-Increment Load&Store operations.
  output logic                      instr_post_incr_valid_o,
  output logic                      lsu_addr_mux_sel_o,
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
  // Signal needed for Hardware Loop operations.
  output logic[31:0] hwlp0_start_o, // To IF stage.
  output logic[31:0] hwlp1_start_o,
//---------------------------------------------------------------------------------



  input  logic                      lsu_addr_incr_req_i,
  input  logic [31:0]               lsu_addr_last_i,



//---------------------------------------------------------------------------------
  // CV-X-IF
  // Issue interface
  output logic                      xif_issue_valid_o,
  output logic [31:0]               xif_issue_req_instr_o,
  input  logic                      xif_issue_ready_i,
  input  logic                      xif_issue_resp_accept_i,
  input  logic                      xif_issue_resp_writeback_i,
  input  logic [2:0]                xif_issue_resp_register_read_i,
  // Register interface
  output logic [31:0]               xif_register_rs1_o,
  output logic [31:0]               xif_register_rs2_o,
  output logic [31:0]               xif_register_rs3_o,
  output logic [2:0]                xif_register_rs_valid_o,
  // Commit interface
  output logic                      xif_commit_valid_o,
  output logic                      xif_commit_kill_o,
  // Result interface
  output logic                      xif_result_ready_o,
  input  logic                      xif_result_valid_i,
  input  logic                      xif_result_we_i,
  input  logic [31:0]               xif_result_data_i,
//---------------------------------------------------------------------------------



  // Interrupt signals
  input  logic                      csr_mstatus_mie_i,
  input  logic                      irq_pending_i,
  input  cve2_pkg::irqs_t           irqs_i,
  input  logic                      irq_nm_i,
  output logic                      nmi_mode_o,

  input  logic                      lsu_load_err_i,
  input  logic                      lsu_store_err_i,

  // Debug Signal
  output logic                      debug_mode_o,
  output cve2_pkg::dbg_cause_e      debug_cause_o,
  output logic                      debug_csr_save_o,
  input  logic                      debug_req_i,
  input  logic                      debug_single_step_i,
  input  logic                      debug_ebreakm_i,
  input  logic                      debug_ebreaku_i,
  input  logic                      trigger_match_i,

  // Write back signal
  input  logic [31:0]               result_ex_i,
  input  logic [31:0]               csr_rdata_i,

  // Register file read
  output logic [4:0]                rf_raddr_a_o,
  input  logic [31:0]               rf_rdata_a_i,
  output logic [4:0]                rf_raddr_b_o,
  input  logic [31:0]               rf_rdata_b_i,



//---------------------------------------------------------------------------------
  output logic [4:0]                rf_raddr_c_o,
  input  logic [31:0]               rf_rdata_c_i,
//---------------------------------------------------------------------------------



  output logic                      rf_ren_a_o,
  output logic                      rf_ren_b_o,



//---------------------------------------------------------------------------------
  output logic                      rf_ren_c_o,
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
  // Register file write (via writeback)
  //1st port.
  output logic [4:0]                rf_waddr_a_id_o,
  output logic [31:0]               rf_wdata_a_id_o,
  output logic                      rf_we_a_id_o,
  //2st port.
  output logic [4:0]                rf_waddr_b_id_o,
  output logic [31:0]               rf_wdata_b_id_o,
  output logic                      rf_we_b_id_o,
//---------------------------------------------------------------------------------



  output  logic                     en_wb_o,
  output  logic                     instr_perf_count_id_o,

  // Performance Counters
  output logic                      perf_jump_o,    // executing a jump instr
  output logic                      perf_branch_o,  // executing a branch instr
  output logic                      perf_tbranch_o, // executing a taken branch instr
  output logic                      perf_dside_wait_o, // instruction in ID/EX is awaiting memory
                                                        // access to finish before proceeding
  output logic                      perf_wfi_wait_o,
  output logic                      perf_div_wait_o,
  output logic                      instr_id_done_o
);

  import cve2_pkg::*;

  // Decoder/Controller, ID stage internal signals
  logic        illegal_insn_dec;
  logic        ebrk_insn;
  logic        mret_insn_dec;
  logic        dret_insn_dec;
  logic        ecall_insn_dec;
  logic        wfi_insn_dec;

  logic        branch_in_dec;
  logic        branch_set, branch_set_raw, branch_set_raw_d;
  logic        branch_jump_set_done_q, branch_jump_set_done_d;
  logic        jump_in_dec;
  logic        jump_set_dec;
  logic        jump_set, jump_set_raw;

  logic        instr_first_cycle;
  logic        instr_executing_spec;
  logic        instr_executing;
  logic        instr_done;
  logic        controller_run;
  logic        stall_mem;
  logic        stall_multdiv;
  logic        stall_branch;
  logic        stall_jump;



//---------------------------------------------------------------------------------
  logic       stall_coproc;
//---------------------------------------------------------------------------------



  logic        stall_id;
  logic        flush_id;
  logic        multicycle_done;

  // Immediate decoding and sign extension
  logic [31:0] imm_i_type;
  logic [31:0] imm_s_type;
  logic [31:0] imm_b_type;
  logic [31:0] imm_u_type;
  logic [31:0] imm_j_type;
  logic [31:0] zimm_rs1_type;



//---------------------------------------------------------------------------------
  logic [31:0] imm_iz_type;
//---------------------------------------------------------------------------------



  logic [31:0] imm_a;       // contains the immediate for operand b
  logic [31:0] imm_b;       // contains the immediate for operand b

  // Register file interface

  rf_wd_sel_e  rf_wdata_sel;
  logic        rf_we_a_dec, rf_we_a_raw;



//---------------------------------------------------------------------------------
  logic        rf_we_b_dec;
//---------------------------------------------------------------------------------



  logic        rf_ren_a, rf_ren_b;



//---------------------------------------------------------------------------------
  logic        rf_ren_c;
//---------------------------------------------------------------------------------



  logic        rf_ren_a_dec, rf_ren_b_dec;



//---------------------------------------------------------------------------------
  logic        rf_ren_c_dec;
//---------------------------------------------------------------------------------



  // Read enables should only be asserted for valid and legal instructions
  assign rf_ren_a = instr_valid_i & ~instr_fetch_err_i & ~illegal_insn_o & rf_ren_a_dec;
  assign rf_ren_b = instr_valid_i & ~instr_fetch_err_i & ~illegal_insn_o & rf_ren_b_dec;



//---------------------------------------------------------------------------------
  assign rf_ren_c = instr_valid_i & ~instr_fetch_err_i & ~illegal_insn_o & rf_ren_c_dec;
//---------------------------------------------------------------------------------



  assign rf_ren_a_o = rf_ren_a;
  assign rf_ren_b_o = rf_ren_b;



//---------------------------------------------------------------------------------
  assign rf_ren_c_o = rf_ren_c;
//---------------------------------------------------------------------------------



  logic [31:0] rf_rdata_a_fwd;
  logic [31:0] rf_rdata_b_fwd;



//---------------------------------------------------------------------------------
  logic [31:0] rf_rdata_c_fwd;
//---------------------------------------------------------------------------------



  // ALU Control
  alu_op_e     alu_operator;
  op_a_sel_e   alu_op_a_mux_sel, alu_op_a_mux_sel_dec;
  op_b_sel_e   alu_op_b_mux_sel, alu_op_b_mux_sel_dec;



//---------------------------------------------------------------------------------
  op_c_sel_e   alu_op_c_mux_sel;
//---------------------------------------------------------------------------------



  logic        alu_multicycle_dec;
  logic        stall_alu;

  logic [33:0] imd_val_q[2];

  imm_a_sel_e  imm_a_mux_sel;
  imm_b_sel_e  imm_b_mux_sel, imm_b_mux_sel_dec;

  // Multiplier Control
  logic        mult_en_id, mult_en_dec; // use integer multiplier
  logic        div_en_id, div_en_dec;   // use integer division or reminder
  logic        multdiv_en_dec;
  md_op_e      multdiv_operator;
  logic [1:0]  multdiv_signed_mode;

  // Data Memory Control
  logic        lsu_we;
  logic [1:0]  lsu_type;
  logic        lsu_sign_ext;
  logic        lsu_req, lsu_req_dec;
  logic        data_req_allowed;

  // CSR control
  logic        csr_pipe_flush;



//---------------------------------------------------------------------------------
 logic        coproc_instr_valid;
 logic        coproc_done;
//---------------------------------------------------------------------------------



  logic [31:0] alu_operand_a;
  logic [31:0] alu_operand_b;



//---------------------------------------------------------------------------------
  logic [31:0] alu_operand_c;
//---------------------------------------------------------------------------------



  /////////////
  // LSU Mux //
  /////////////

  // Misaligned loads/stores result in two aligned loads/stores, compute second address
  assign alu_op_a_mux_sel = lsu_addr_incr_req_i ? OP_A_FWD        : alu_op_a_mux_sel_dec;
  assign alu_op_b_mux_sel = lsu_addr_incr_req_i ? OP_B_IMM        : alu_op_b_mux_sel_dec;
  assign imm_b_mux_sel    = lsu_addr_incr_req_i ? IMM_B_INCR_ADDR : imm_b_mux_sel_dec;

  ///////////////////
  // Operand MUXES //
  ///////////////////

  // Main ALU immediate MUX for Operand A
  assign imm_a = (imm_a_mux_sel == IMM_A_Z) ? zimm_rs1_type : '0;

  // Main ALU MUX for Operand A
  always_comb begin : alu_operand_a_mux
    unique case (alu_op_a_mux_sel)
      OP_A_REG_A:  alu_operand_a = rf_rdata_a_fwd;
      OP_A_FWD:    alu_operand_a = lsu_addr_last_i;
      OP_A_CURRPC: alu_operand_a = pc_id_i;
      OP_A_IMM:    alu_operand_a = imm_a;
      default:     alu_operand_a = pc_id_i;
    endcase
  end

  op_a_sel_e  unused_a_mux_sel;
  imm_b_sel_e unused_b_mux_sel;

  // Full main ALU immediate MUX for Operand B
  always_comb begin : immediate_b_mux
    unique case (imm_b_mux_sel)
      IMM_B_I:         imm_b = imm_i_type;
      IMM_B_S:         imm_b = imm_s_type;
      IMM_B_B:         imm_b = imm_b_type;
      IMM_B_U:         imm_b = imm_u_type;
      IMM_B_J:         imm_b = imm_j_type;
      IMM_B_INCR_PC:   imm_b = instr_is_compressed_i ? 32'h2 : 32'h4;
      IMM_B_INCR_ADDR: imm_b = 32'h4;
      default:         imm_b = 32'h4;
    endcase
  end
  `ASSERT(IbexImmBMuxSelValid, instr_valid_i |-> imm_b_mux_sel inside {
      IMM_B_I,
      IMM_B_S,
      IMM_B_B,
      IMM_B_U,
      IMM_B_J,
      IMM_B_INCR_PC,
      IMM_B_INCR_ADDR})



//---------------------------------------------------------------------------------
  // Operand C MUX: needed for Register-Register Stores with Post-Increment and Register-Register Stores.
  // The adder needs rs1 and rs3 as inputs to calculate the incremented address (Register-Register Stores with Post-Increment: rs1+=rs3) 
  // or to calculate the actual adress (Register-Register Stores: Mem(rs1+rs3)). Therefore, rs3 is routed by means of the MUX for Operand B 
  // to the second input of the adder whereas the data to be stored pass through ALU Operand C.

  always_comb begin : alu_operand_b_mux
    unique case (alu_op_b_mux_sel)
      OP_B_REG_B: alu_operand_b = rf_rdata_b_fwd;
      OP_B_IMM:   alu_operand_b = imm_b;
      OP_B_REG_C: alu_operand_b = rf_rdata_c_fwd;
    endcase
  end

  always_comb begin : alu_operand_c_mux
    unique case (alu_op_c_mux_sel)
      OP_C_REG_C:  alu_operand_c = rf_rdata_c_fwd;
      OP_C_REG_B:  alu_operand_c = rf_rdata_b_fwd;
    endcase
  end
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
  // Hardware Loop.

  // Intermediate signals,
  // hwloop_regs input signals.
  logic [1:0]               hwlp_start_mux_sel;
  logic [31:0]              hwlp_start_d;
  logic [1:0]               hwlp_end_mux_sel;
  logic [31:0]              hwlp_end_d;
  logic                     hwlp_cnt_mux_sel;
  logic [31:0]              hwlp_cnt_d;
  logic [2:0]               hwlp_we;
  logic                     hwlp_regid;

  // hwloops_regs output signals.
  logic [N_HWLP-1:0][31:0]  hwlp_start_q; // To IF stage.
  logic [N_HWLP-1:0][31:0]  hwlp_end_q;   // To controller.
  logic [N_HWLP-1:0][31:0]  hwlp_cnt_q;   // 

  assign hwlp0_start_o = hwlp_start_q[0];
  assign hwlp1_start_o = hwlp_start_q[1];

  // Counter enable (from controller to hwloop_regs)
  logic[N_HWLP-1:0]         hwlp_dec_cnt; 

  //Start address.
  always_comb begin
    case (hwlp_start_mux_sel)
      2'b00:   hwlp_start_d = hwlp_end_d;  
      2'b01:   hwlp_start_d = pc_id_i + 4;  
      2'b10:   hwlp_start_d = rf_rdata_a_fwd;
      default: hwlp_start_d = rf_rdata_a_fwd;
    endcase
  end

  //End address.
  always_comb begin
    case (hwlp_end_mux_sel)
      2'b00:   hwlp_end_d = pc_id_i + {imm_iz_type[29:0], 2'b0};
      2'b01:   hwlp_end_d = pc_id_i + {zimm_rs1_type[29:0], 2'b0};
      2'b10:   hwlp_end_d = rf_rdata_a_fwd;
      default: hwlp_end_d = rf_rdata_a_fwd;
    endcase
  end

  //Counter value.
  always_comb begin : hwlp_cnt_mux
    case (hwlp_cnt_mux_sel)
      1'b0: hwlp_cnt_d = imm_iz_type;
      1'b1: hwlp_cnt_d = rf_rdata_a_fwd;
    endcase
    ;
  end

  assign hwlp_regid = instr_rdata_i[7];

  cve2_hwloop_regs #(
    .N_REGS(N_HWLP)
  )
  cve2_hwloop_regs_i (
    .clk(clk_i),
    .rst_n(rst_ni),


    .hwlp_start_data_i(hwlp_start_d),
    .hwlp_end_data_i  (hwlp_end_d),
    .hwlp_cnt_data_i  (hwlp_cnt_d),
    .hwlp_we_i        (hwlp_we),
    .hwlp_regid_i     (hwlp_regid),  


    .valid_i(instr_valid_i),


    .hwlp_dec_cnt_i(hwlp_dec_cnt), 


    .hwlp_start_addr_o(hwlp_start_q),
    .hwlp_end_addr_o  (hwlp_end_q),
    .hwlp_counter_o   (hwlp_cnt_q)
  );

//---------------------------------------------------------------------------------



  /////////////////////////////////////////
  // Multicycle Operation Stage Register //
  /////////////////////////////////////////

  for (genvar i = 0; i < 2; i++) begin : gen_intermediate_val_reg
    always_ff @(posedge clk_i or negedge rst_ni) begin : intermediate_val_reg
      if (!rst_ni) begin
        imd_val_q[i] <= '0;
      end else if (imd_val_we_ex_i[i]) begin
        imd_val_q[i] <= imd_val_d_ex_i[i];
      end
    end
  end

  assign imd_val_q_ex_o = imd_val_q;

  ///////////////////////
  // Register File MUX //
  ///////////////////////

  // Suppress register write if there is an illegal CSR access or instruction is not executing
  assign rf_we_a_id_o = rf_we_a_raw & instr_executing & ~illegal_csr_insn_i;



//---------------------------------------------------------------------------------
  //The 2nd register file write port is not involved in CSR operations.
  assign rf_we_b_id_o =  rf_we_b_dec & instr_executing;
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
  // 1st register file write port data mux.
  always_comb begin : rf_wdata_id_mux
    unique case (rf_wdata_sel)
      RF_WD_EX:     rf_wdata_a_id_o = result_ex_i;
      RF_WD_CSR:    rf_wdata_a_id_o = csr_rdata_i;
      RF_WD_COPROC: rf_wdata_a_id_o = xif_result_data_i;
      default:      rf_wdata_a_id_o = result_ex_i;
    endcase
  end

  // 2nd register file write port data.
  assign rf_wdata_b_id_o = result_ex_i;
//---------------------------------------------------------------------------------



  /////////////
  // Decoder //
  /////////////

  cve2_decoder #(
    .RV32E          (RV32E),
    .RV32M          (RV32M),
    .RV32B          (RV32B),
    .COPROC_OPCODE  (COPROC_OPCODE)
  ) decoder_i (
    .clk_i (clk_i),
    .rst_ni(rst_ni),
    // controller
    .illegal_insn_o(illegal_insn_dec),
    .ebrk_insn_o   (ebrk_insn),
    .mret_insn_o   (mret_insn_dec),
    .dret_insn_o   (dret_insn_dec),
    .ecall_insn_o  (ecall_insn_dec),
    .wfi_insn_o    (wfi_insn_dec),
    .jump_set_o    (jump_set_dec),

    // from IF-ID pipeline register
    .instr_first_cycle_i(instr_first_cycle),
    .instr_rdata_i      (instr_rdata_i),
    .instr_rdata_alu_i  (instr_rdata_alu_i),
    .illegal_c_insn_i   (illegal_c_insn_i),

    // immediates
    .imm_a_mux_sel_o(imm_a_mux_sel),
    .imm_b_mux_sel_o(imm_b_mux_sel_dec),

    .imm_i_type_o   (imm_i_type),
    .imm_s_type_o   (imm_s_type),
    .imm_b_type_o   (imm_b_type),
    .imm_u_type_o   (imm_u_type),
    .imm_j_type_o   (imm_j_type),
    .zimm_rs1_type_o(zimm_rs1_type),
    .imm_iz_type_o  (imm_iz_type),

    // register file
    .rf_wdata_sel_o(rf_wdata_sel),
    .rf_we_a_o     (rf_we_a_dec),



//---------------------------------------------------------------------------------
    .rf_we_b_o(rf_we_b_dec),
//---------------------------------------------------------------------------------



    .rf_raddr_a_o(rf_raddr_a_o),
    .rf_raddr_b_o(rf_raddr_b_o),



//---------------------------------------------------------------------------------
    .rf_raddr_c_o(rf_raddr_c_o),
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
    .rf_waddr_a_o(rf_waddr_a_id_o),
    .rf_waddr_b_o(rf_waddr_b_id_o),
//---------------------------------------------------------------------------------



    .rf_ren_a_o  (rf_ren_a_dec),
    .rf_ren_b_o  (rf_ren_b_dec),



//---------------------------------------------------------------------------------
    .rf_ren_c_o  (rf_ren_c_dec),
//---------------------------------------------------------------------------------



    // ALU
    .alu_operator_o    (alu_operator),
    .alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),



//---------------------------------------------------------------------------------
    .alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
    .alu_op_c_mux_sel_o(alu_op_c_mux_sel),    
//---------------------------------------------------------------------------------



    .alu_multicycle_o  (alu_multicycle_dec),

    // MULT & DIV
    .mult_en_o            (mult_en_dec),
    .div_en_o             (div_en_dec),
    .mult_sel_o           (mult_sel_ex_o),
    .div_sel_o            (div_sel_ex_o),
    .multdiv_operator_o   (multdiv_operator),
    .multdiv_signed_mode_o(multdiv_signed_mode),

    // CSRs
    .csr_access_o(csr_access_o),
    .csr_op_o    (csr_op_o),

    // LSU
    .data_req_o           (lsu_req_dec),
    .data_we_o            (lsu_we),
    .data_type_o          (lsu_type),
    .data_sign_extension_o(lsu_sign_ext),



//---------------------------------------------------------------------------------
    .hwlp_start_mux_sel_o(hwlp_start_mux_sel), 
    .hwlp_end_mux_sel_o  (hwlp_end_mux_sel),   
    .hwlp_cnt_mux_sel_o  (hwlp_cnt_mux_sel),   
    .hwlp_we_o           (hwlp_we),            
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
    .instr_post_incr_valid_o(instr_post_incr_valid_o),
    .lsu_addr_mux_sel_o(lsu_addr_mux_sel_o), 
//---------------------------------------------------------------------------------



//---------------------------------------------------------------------------------
    .xif_issue_resp_register_read_i(xif_issue_resp_register_read_i),
    .xif_issue_resp_writeback_i(xif_issue_resp_writeback_i),
    .coproc_instr_valid_o(coproc_instr_valid),
//---------------------------------------------------------------------------------





    // jump/branches
    .jump_in_dec_o  (jump_in_dec),
    .branch_in_dec_o(branch_in_dec)
  );

  /////////////////////////////////
  // CSR-related pipeline flushes //
  /////////////////////////////////
  always_comb begin : csr_pipeline_flushes
    csr_pipe_flush = 1'b0;

    // A pipeline flush is needed to let the controller react after modifying certain CSRs:
    // - When enabling interrupts, pending IRQs become visible to the controller only during
    //   the next cycle. If during that cycle the core disables interrupts again, it does not
    //   see any pending IRQs and consequently does not start to handle interrupts.
    // - When modifying any PMP CSR, PMP check of the next instruction might get invalidated.
    //   Hence, a pipeline flush is needed to instantiate another PMP check with the updated CSRs.
    // - When modifying debug CSRs - TODO: Check if this is really needed
    if (csr_op_en_o == 1'b1 && (csr_op_o == CSR_OP_WRITE || csr_op_o == CSR_OP_SET)) begin
      if (csr_num_e'(instr_rdata_i[31:20]) == CSR_MSTATUS ||
          csr_num_e'(instr_rdata_i[31:20]) == CSR_MIE     ||
          csr_num_e'(instr_rdata_i[31:20]) == CSR_MSECCFG ||
          // To catch all PMPCFG/PMPADDR registers, get the shared top most 7 bits.
          instr_rdata_i[31:25] == 7'h1D) begin
        csr_pipe_flush = 1'b1;
      end
    end else if (csr_op_en_o == 1'b1 && csr_op_o != CSR_OP_READ) begin
      if (csr_num_e'(instr_rdata_i[31:20]) == CSR_DCSR      ||
          csr_num_e'(instr_rdata_i[31:20]) == CSR_DPC       ||
          csr_num_e'(instr_rdata_i[31:20]) == CSR_DSCRATCH0 ||
          csr_num_e'(instr_rdata_i[31:20]) == CSR_DSCRATCH1) begin
        csr_pipe_flush = 1'b1;
      end
    end
  end

  ////////////////
  // Controller //
  ////////////////

//---------------------------------------------------------------------------------
  assign illegal_insn_o = instr_valid_i && (illegal_insn_dec || illegal_csr_insn_i || (xif_issue_valid_o && xif_issue_ready_i && ~xif_issue_resp_accept_i));
//---------------------------------------------------------------------------------

  cve2_controller #(
    .N_HWLP      (N_HWLP)
  ) controller_i (
    .clk_i (clk_i),
    .rst_ni(rst_ni),

    .fetch_enable_i(fetch_enable_i),
    .ctrl_busy_o(ctrl_busy_o),

    // decoder related signals
    .illegal_insn_i  (illegal_insn_o),
    .ecall_insn_i    (ecall_insn_dec),
    .mret_insn_i     (mret_insn_dec),
    .dret_insn_i     (dret_insn_dec),
    .wfi_insn_i      (wfi_insn_dec),
    .ebrk_insn_i     (ebrk_insn),
    .csr_pipe_flush_i(csr_pipe_flush),

    // from IF-ID pipeline
    .instr_valid_i          (instr_valid_i),
    .instr_i                (instr_rdata_i),
    .instr_compressed_i     (instr_rdata_c_i),
    .instr_is_compressed_i  (instr_is_compressed_i),
    .instr_fetch_err_i      (instr_fetch_err_i),
    .instr_fetch_err_plus2_i(instr_fetch_err_plus2_i),
    .pc_id_i                (pc_id_i),

    // to IF-ID pipeline
    .instr_valid_clear_o(instr_valid_clear_o),
    .id_in_ready_o      (id_in_ready_o),
    .controller_run_o   (controller_run),

    // to prefetcher
    .instr_req_o           (instr_req_o),
    .pc_set_o              (pc_set_o),
    .pc_mux_o              (pc_mux_o),
    .exc_pc_mux_o          (exc_pc_mux_o),
    .exc_cause_o           (exc_cause_o),

    // LSU
    .lsu_addr_last_i(lsu_addr_last_i),
    .load_err_i     (lsu_load_err_i),
    .store_err_i    (lsu_store_err_i),
    // jump/branch control
    .branch_set_i     (branch_set),
    .jump_set_i       (jump_set),

    // interrupt signals
    .csr_mstatus_mie_i(csr_mstatus_mie_i),
    .irq_pending_i    (irq_pending_i),
    .irqs_i           (irqs_i),
    .irq_nm_i         (irq_nm_i),
    .nmi_mode_o       (nmi_mode_o),

    // CSR Controller Signals
    .csr_save_if_o        (csr_save_if_o),
    .csr_save_id_o        (csr_save_id_o),
    .csr_restore_mret_id_o(csr_restore_mret_id_o),
    .csr_restore_dret_id_o(csr_restore_dret_id_o),
    .csr_save_cause_o     (csr_save_cause_o),
    .csr_mtval_o          (csr_mtval_o),
    .priv_mode_i          (priv_mode_i),
    .csr_mstatus_tw_i     (csr_mstatus_tw_i),

    // Debug Signal
    .debug_mode_o       (debug_mode_o),
    .debug_cause_o      (debug_cause_o),
    .debug_csr_save_o   (debug_csr_save_o),
    .debug_req_i        (debug_req_i),
    .debug_single_step_i(debug_single_step_i),
    .debug_ebreakm_i    (debug_ebreakm_i),
    .debug_ebreaku_i    (debug_ebreaku_i),
    .trigger_match_i    (trigger_match_i),

    .stall_id_i(stall_id),
    .flush_id_o(flush_id),

    // Performance Counters
    .perf_jump_o   (perf_jump_o),
    .perf_tbranch_o(perf_tbranch_o),



  //---------------------------------------------------------------------------------
    .hwlp_end_i(hwlp_start_q),
    .hwlp_cnt_i(hwlp_cnt_q),
    .hwlp_dec_cnt_o(hwlp_dec_cnt)
  //---------------------------------------------------------------------------------


  
  );

  assign multdiv_en_dec   = mult_en_dec | div_en_dec;

  assign lsu_req         = instr_executing ? data_req_allowed & lsu_req_dec  : 1'b0;
  assign mult_en_id      = instr_executing ? mult_en_dec                     : 1'b0;
  assign div_en_id       = instr_executing ? div_en_dec                      : 1'b0;

  assign lsu_req_o               = lsu_req;
  assign lsu_we_o                = lsu_we;
  assign lsu_type_o              = lsu_type;
  assign lsu_sign_ext_o          = lsu_sign_ext;
  assign lsu_wdata_o             = rf_rdata_b_fwd;
  // csr_op_en_o is set when CSR access should actually happen.
  // csv_access_o is set when CSR access instruction is present and is used to compute whether a CSR
  // access is illegal. A combinational loop would be created if csr_op_en_o was used along (as
  // asserting it for an illegal csr access would result in a flush that would need to deassert it).
  assign csr_op_en_o             = csr_access_o & instr_executing & instr_id_done_o;

  assign alu_operator_ex_o           = alu_operator;
  assign alu_operand_a_ex_o          = alu_operand_a;
  assign alu_operand_b_ex_o          = alu_operand_b;



//---------------------------------------------------------------------------------
  assign alu_operand_c_ex_o          = alu_operand_c;
//---------------------------------------------------------------------------------



  assign mult_en_ex_o                = mult_en_id;
  assign div_en_ex_o                 = div_en_id;

  assign multdiv_operator_ex_o       = multdiv_operator;
  assign multdiv_signed_mode_ex_o    = multdiv_signed_mode;
  assign multdiv_operand_a_ex_o      = rf_rdata_a_fwd;
  assign multdiv_operand_b_ex_o      = rf_rdata_b_fwd;



//---------------------------------------------------------------------------------
  assign xif_issue_req_instr_o       = instr_rdata_i;
  assign xif_register_rs1_o          = rf_rdata_a_fwd;
  assign xif_register_rs2_o          = rf_rdata_b_fwd;
  assign xif_register_rs3_o          = rf_rdata_c_fwd; 

  logic commit_valid_q, commit_valid_d;
  assign commit_valid_d = xif_issue_valid_o && xif_issue_ready_i && xif_issue_resp_accept_i;
  always_ff@(posedge clk_i or negedge rst_ni) begin
    if(~rst_ni) begin
      commit_valid_q <= 1'b0;
    end
    else begin
      commit_valid_q <= commit_valid_d;
    end
  end

  assign xif_commit_valid_o = commit_valid_q;

  assign xif_commit_kill_o = 1'b0;
  
  assign xif_result_ready_o = 1'b1;
//---------------------------------------------------------------------------------



  ////////////////////////
  // Branch set control //
  ////////////////////////

  // SEC_CM: CORE.DATA_REG_SW.SCA
  // Branch set flopped without branch target ALU, or in fixed time execution mode
  // (condition pass/fail used next cycle where branch target is calculated)
  logic branch_set_raw_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      branch_set_raw_q <= 1'b0;
    end else begin
      branch_set_raw_q <= branch_set_raw_d;
    end
  end

  // Branches always take two cycles in fixed time execution mode, with or without the branch
  // target ALU (to avoid a path from the branch decision into the branch target ALU operand
  // muxing).
  assign branch_set_raw      = branch_set_raw_q;


  // Track whether the current instruction in ID/EX has done a branch or jump set.
  assign branch_jump_set_done_d = (branch_set_raw | jump_set_raw | branch_jump_set_done_q) &
    ~instr_valid_clear_o;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      branch_jump_set_done_q <= 1'b0;
    end else begin
      branch_jump_set_done_q <= branch_jump_set_done_d;
    end
  end

  // the _raw signals from the state machine may be asserted for multiple cycles when
  // instr_executing_spec is asserted and instr_executing is not asserted. This may occur where
  // a memory error is seen or a there are outstanding memory accesses (indicate a load or store is
  // in the WB stage). The branch or jump speculatively begins the fetch but is held back from
  // completing until it is certain the outstanding access hasn't seen a memory error. This logic
  // ensures only the first cycle of a branch or jump set is sent to the controller to prevent
  // needless extra IF flushes and fetches.
  assign jump_set        = jump_set_raw        & ~branch_jump_set_done_q;
  assign branch_set      = branch_set_raw      & ~branch_jump_set_done_q;

  ///////////////
  // ID-EX FSM //
  ///////////////

  typedef enum logic { FIRST_CYCLE, MULTI_CYCLE } id_fsm_e;
  id_fsm_e id_fsm_q, id_fsm_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin : id_pipeline_reg
    if (!rst_ni) begin
      id_fsm_q <= FIRST_CYCLE;
    end else if (instr_executing) begin
      id_fsm_q <= id_fsm_d;
    end
  end

  // ID/EX stage can be in two states, FIRST_CYCLE and MULTI_CYCLE. An instruction enters
  // MULTI_CYCLE if it requires multiple cycles to complete regardless of stalls and other
  // considerations. An instruction may be held in FIRST_CYCLE if it's unable to begin executing
  // (this is controlled by instr_executing).

  always_comb begin
    id_fsm_d                = id_fsm_q;
    rf_we_a_raw             = rf_we_a_dec;
    stall_multdiv           = 1'b0;
    stall_jump              = 1'b0;
    stall_branch            = 1'b0;
    stall_alu               = 1'b0;

  //---------------------------------------------------------------------------------
    //xif_commit_valid_o    = 1'b0;
    stall_coproc            = 1'b0;
  //---------------------------------------------------------------------------------

    branch_set_raw_d        = 1'b0;
    jump_set_raw            = 1'b0;
    perf_branch_o           = 1'b0;

    if (instr_executing_spec) begin
      unique case (id_fsm_q)
        FIRST_CYCLE: begin
          unique case (1'b1)
            lsu_req_dec: begin
              begin
                // LSU operation
                id_fsm_d    = MULTI_CYCLE;
              end
            end
            multdiv_en_dec: begin
              // MUL or DIV operation
              if (~ex_valid_i) begin
                // When single-cycle multiply is configured mul can finish in the first cycle so
                // only enter MULTI_CYCLE state if a result isn't immediately available
                id_fsm_d      = MULTI_CYCLE;
                rf_we_a_raw   = 1'b0;
                stall_multdiv = 1'b1;
              end
            end
            branch_in_dec: begin
              // cond branch operation
              // All branches take two cycles in fixed time execution mode, regardless of branch
              // condition.
              // SEC_CM: CORE.DATA_REG_SW.SCA
              id_fsm_d         = (branch_decision_i) ?
                                     MULTI_CYCLE : FIRST_CYCLE;
              stall_branch     = branch_decision_i;
              branch_set_raw_d = branch_decision_i;

              perf_branch_o = 1'b1;
            end
            jump_in_dec: begin
              // uncond branch operation
              id_fsm_d      = MULTI_CYCLE;
              stall_jump    = 1'b1;
              jump_set_raw  = jump_set_dec;
            end
            alu_multicycle_dec: begin
              stall_alu     = 1'b1;
              id_fsm_d      = MULTI_CYCLE;
              rf_we_a_raw   = 1'b0;
            end

//---------------------------------------------------------------------------------
            coproc_instr_valid: begin
              if (xif_issue_ready_i && xif_issue_resp_writeback_i) begin
                id_fsm_d             = MULTI_CYCLE;
                //xif_commit_valid_o = 1'b1;
              end
              stall_coproc = ~xif_issue_ready_i || xif_issue_resp_writeback_i; 
              rf_we_a_raw  = 1'b0;
            end
//---------------------------------------------------------------------------------

            default: begin
              id_fsm_d      = FIRST_CYCLE;
            end
          endcase
        end

        MULTI_CYCLE: begin
          if(multdiv_en_dec) begin
            rf_we_a_raw       = rf_we_a_dec & ex_valid_i;
          end

          if (multicycle_done) begin
            id_fsm_d        = FIRST_CYCLE;
          end else begin
            stall_multdiv   = multdiv_en_dec;
            stall_branch    = branch_in_dec;
            stall_jump      = jump_in_dec;

//---------------------------------------------------------------------------------
            stall_coproc    = coproc_instr_valid;
//---------------------------------------------------------------------------------

          end
        end

        default: begin
          id_fsm_d          = FIRST_CYCLE;
        end
      endcase
    end
  end

//---------------------------------------------------------------------------------  
  assign xif_issue_valid_o = instr_executing && coproc_instr_valid && (id_fsm_q == FIRST_CYCLE);
  assign coproc_done       = (xif_issue_valid_o && xif_issue_ready_i && ~xif_issue_resp_writeback_i) || (xif_result_valid_i && xif_result_we_i);
//---------------------------------------------------------------------------------

  `ASSERT(StallIDIfMulticycle, (id_fsm_q == FIRST_CYCLE) & (id_fsm_d == MULTI_CYCLE) |-> stall_id)


  // Stall ID/EX stage for reason that relates to instruction in ID/EX, update assertion below if
  // modifying this.

//---------------------------------------------------------------------------------
  assign stall_id = stall_mem | stall_multdiv | stall_jump | stall_branch |
                      stall_alu | stall_coproc;
//---------------------------------------------------------------------------------

  // Generally illegal instructions have no reason to stall, however they must still stall waiting
  // for outstanding memory requests so exceptions related to them take priority over the illegal
  // instruction exception.
  `ASSERT(IllegalInsnStallMustBeMemStall, illegal_insn_o & stall_id |-> stall_mem &
    ~(stall_multdiv | stall_jump | stall_branch | stall_alu))

  assign instr_done = ~stall_id & ~flush_id & instr_executing;

  // Signal instruction in ID is in it's first cycle. It can remain in its
  // first cycle if it is stalled.
  assign instr_first_cycle      = instr_valid_i & (id_fsm_q == FIRST_CYCLE);
  // Used by RVFI to know when to capture register read data
  // Used by ALU to access RS3 if ternary instruction.
  assign instr_first_cycle_id_o = instr_first_cycle;

    assign multicycle_done = lsu_req_dec ? lsu_resp_valid_i :
                             (coproc_instr_valid ? coproc_done : ex_valid_i);

    assign data_req_allowed = instr_first_cycle;

    // Without Writeback Stage always stall the first cycle of a load/store.
    // Then stall until it is complete
    assign stall_mem = instr_valid_i & (lsu_req_dec & (~lsu_resp_valid_i | instr_first_cycle));

    // Without writeback stage any valid instruction that hasn't seen an error will execute
    assign instr_executing_spec = instr_valid_i & ~instr_fetch_err_i & controller_run;
    assign instr_executing = instr_executing_spec;

    `ASSERT(IbexStallIfValidInstrNotExecuting,
      instr_valid_i & ~instr_fetch_err_i & ~instr_executing & controller_run |-> stall_id)

    // No data forwarding without writeback stage so always take source register data direct from
    // register file
    assign rf_rdata_a_fwd = rf_rdata_a_i;
    assign rf_rdata_b_fwd = rf_rdata_b_i;

//---------------------------------------------------------------------------------
    assign rf_rdata_c_fwd  = rf_rdata_c_i;
//---------------------------------------------------------------------------------

//---------------------------------------------------------------------------------
    //Since hazard can not occour all the source registers are always valid.
    assign xif_register_rs_valid_o[0] = 1'b1;
    assign xif_register_rs_valid_o[1] = 1'b1;
    assign xif_register_rs_valid_o[2] = 1'b1;
//--------------------------------------------------------------------------------- 

    // Unused Writeback stage only IO & wiring
    // Assign inputs and internal wiring to unused signals to satisfy lint checks
    // Tie-off outputs to constant values
    logic unused_data_req_done_ex;

    assign perf_dside_wait_o = instr_executing & lsu_req_dec & ~lsu_resp_valid_i;

    assign instr_id_done_o = instr_done;

  // Signal which instructions to count as retired in minstret, all traps along with ebrk and
  // ecall instructions are not counted.
  assign instr_perf_count_id_o = ~ebrk_insn & ~ecall_insn_dec & ~illegal_insn_dec &
      ~(dret_insn_dec & ~debug_mode_o) &
      ~illegal_csr_insn_i & ~instr_fetch_err_i;

  // An instruction is ready to move to the writeback
  assign en_wb_o = instr_done;

  assign perf_wfi_wait_o = wfi_insn_dec;
  assign perf_div_wait_o = stall_multdiv & div_en_dec;

  //////////
  // FCOV //
  //////////

  `DV_FCOV_SIGNAL(logic, branch_taken,
    instr_executing & (id_fsm_q == FIRST_CYCLE) & branch_decision_i)
  `DV_FCOV_SIGNAL(logic, branch_not_taken,
    instr_executing & (id_fsm_q == FIRST_CYCLE) & ~branch_decision_i)

  ////////////////
  // Assertions //
  ////////////////

  // Selectors must be known/valid.
  `ASSERT_KNOWN_IF(IbexAluOpMuxSelKnown, alu_op_a_mux_sel, instr_valid_i)
  `ASSERT(IbexAluAOpMuxSelValid, instr_valid_i |-> alu_op_a_mux_sel inside {
      OP_A_REG_A,
      OP_A_FWD,
      OP_A_CURRPC,
      OP_A_IMM})
  `ASSERT(IbexRegfileWdataSelValid, instr_valid_i |-> rf_wdata_sel inside {
      RF_WD_EX,
      RF_WD_CSR, 
      RF_WD_COPROC})
  `ASSERT_KNOWN(IbexWbStateKnown, id_fsm_q)

  // Branch decision must be valid when jumping.
  `ASSERT_KNOWN_IF(IbexBranchDecisionValid, branch_decision_i,
      instr_valid_i && !(illegal_csr_insn_i || instr_fetch_err_i))

  // Instruction delivered to ID stage can not contain X.
  `ASSERT_KNOWN_IF(IbexIdInstrKnown, instr_rdata_i,
      instr_valid_i && !(illegal_c_insn_i || instr_fetch_err_i))

  // Instruction delivered to ID stage can not contain X.
  `ASSERT_KNOWN_IF(IbexIdInstrALUKnown, instr_rdata_alu_i,
      instr_valid_i && !(illegal_c_insn_i || instr_fetch_err_i))

  // Multicycle enable signals must be unique.
  `ASSERT(IbexMulticycleEnableUnique,
      $onehot0({lsu_req_dec, multdiv_en_dec, branch_in_dec, jump_in_dec}))

  // Duplicated instruction flops must match
  // === as DV environment can produce instructions with Xs in, so must use precise match that
  // includes Xs
  `ASSERT(IbexDuplicateInstrMatch, instr_valid_i |-> instr_rdata_i === instr_rdata_alu_i)

  `ifdef CHECK_MISALIGNED
  `ASSERT(IbexMisalignedMemoryAccess, !lsu_addr_incr_req_i)
  `endif

endmodule
